module Alu ();

endmodule
